module two_state();

real       pi;
bit [3:0] bit_test; 
byte      byte_test; // same as above
initial begin
   pi             = 3.1415;
   bit_test       = 4'd7;
   byte_test      = 4'd7;
end

endmodule